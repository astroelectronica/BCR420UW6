.title KiCad schematic
.include "C:/AE/BCR420UW6/BCR420UW6.spice.txt"
.include "C:/AE/BCR420UW6/SML-011VT_SPICE.lib"
D2 /LD1 /LD2 SML-011VT
D3 /LD2 /LD3 SML-011VT
D1 VCC /LD1 SML-011VT
XU1 /EN /LD4 /LD4 0 /LD4 /REXT BCR420UW6
D4 /LD3 /LD4 SML-011VT
V1 VCC 0 DC {VSOURCE} 
R1 /REXT 0 {REXT}
V2 /EN 0 DC {EN} 
.end
